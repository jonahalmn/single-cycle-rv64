module debug_gpr #(parameter ARCH_WIDTH = 64) (input wire[31:0][ARCH_WIDTH - 1:0]regsData);

wire[ARCH_WIDTH - 1:0] zero;
wire[ARCH_WIDTH - 1:0] ra;
wire[ARCH_WIDTH - 1:0] sp;
wire[ARCH_WIDTH - 1:0] gp;
wire[ARCH_WIDTH - 1:0] tp;
wire[ARCH_WIDTH - 1:0] t0;
wire[ARCH_WIDTH - 1:0] t1;
wire[ARCH_WIDTH - 1:0] t2;
wire[ARCH_WIDTH - 1:0] s0;
wire[ARCH_WIDTH - 1:0] s1;
wire[ARCH_WIDTH - 1:0] a0;
wire[ARCH_WIDTH - 1:0] a1;
wire[ARCH_WIDTH - 1:0] a2;
wire[ARCH_WIDTH - 1:0] a3;
wire[ARCH_WIDTH - 1:0] a4;
wire[ARCH_WIDTH - 1:0] a5;
wire[ARCH_WIDTH - 1:0] a6;
wire[ARCH_WIDTH - 1:0] a7;
wire[ARCH_WIDTH - 1:0] s2;
wire[ARCH_WIDTH - 1:0] s3;
wire[ARCH_WIDTH - 1:0] s4;
wire[ARCH_WIDTH - 1:0] s5;
wire[ARCH_WIDTH - 1:0] s6;
wire[ARCH_WIDTH - 1:0] s7;
wire[ARCH_WIDTH - 1:0] s8;
wire[ARCH_WIDTH - 1:0] s9;
wire[ARCH_WIDTH - 1:0] s10;
wire[ARCH_WIDTH - 1:0] s11;
wire[ARCH_WIDTH - 1:0] t3;
wire[ARCH_WIDTH - 1:0] t4;
wire[ARCH_WIDTH - 1:0] t5;
wire[ARCH_WIDTH - 1:0] t6;

assign zero = regsData[0];
assign ra = regsData[1];
assign sp = regsData[2];
assign gp = regsData[3];
assign tp = regsData[4];
assign t0 = regsData[5];
assign t1 = regsData[6];
assign t2 = regsData[7];
assign s0 = regsData[8];
assign s1 = regsData[9];
assign a0 = regsData[10];
assign a1 = regsData[11];
assign a2 = regsData[12];
assign a3 = regsData[13];
assign a4 = regsData[14];
assign a5 = regsData[15];
assign a6 = regsData[16];
assign a7 = regsData[17];
assign s2 = regsData[18];
assign s3 = regsData[19];
assign s4 = regsData[20];
assign s5 = regsData[21];
assign s6 = regsData[22];
assign s7 = regsData[23];
assign s8 = regsData[24];
assign s9 = regsData[25];
assign s10 = regsData[26];
assign s11 = regsData[27];
assign t3 = regsData[28];
assign t4 = regsData[29];
assign t5 = regsData[30];
assign t6 = regsData[31];

endmodule